// final_soc.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module final_soc (
		input  wire          clk_clk,                //             clk.clk
		input  wire          frame_sync_export,      //      frame_sync.export
		output wire [2047:0] gamefile_export_data,   //        gamefile.export_data
		output wire [1:0]    otg_hpi_address_export, // otg_hpi_address.export
		output wire          otg_hpi_cs_export,      //      otg_hpi_cs.export
		input  wire [15:0]   otg_hpi_data_in_port,   //    otg_hpi_data.in_port
		output wire [15:0]   otg_hpi_data_out_port,  //                .out_port
		output wire          otg_hpi_r_export,       //       otg_hpi_r.export
		output wire          otg_hpi_reset_export,   //   otg_hpi_reset.export
		output wire          otg_hpi_w_export,       //       otg_hpi_w.export
		input  wire          reset_reset_n,          //           reset.reset_n
		output wire          sdram_clk_clk,          //       sdram_clk.clk
		output wire [12:0]   sdram_wire_addr,        //      sdram_wire.addr
		output wire [1:0]    sdram_wire_ba,          //                .ba
		output wire          sdram_wire_cas_n,       //                .cas_n
		output wire          sdram_wire_cke,         //                .cke
		output wire          sdram_wire_cs_n,        //                .cs_n
		inout  wire [31:0]   sdram_wire_dq,          //                .dq
		output wire [3:0]    sdram_wire_dqm,         //                .dqm
		output wire          sdram_wire_ras_n,       //                .ras_n
		output wire          sdram_wire_we_n         //                .we_n
	);

	wire         system_pll_c0_clk;                                         // system_pll:c0 -> [mm_interconnect_0:system_pll_c0_clk, rst_controller_002:clk, sdram:clk]
	wire  [31:0] game_cpu_data_master_readdata;                             // mm_interconnect_0:game_cpu_data_master_readdata -> game_cpu:d_readdata
	wire         game_cpu_data_master_waitrequest;                          // mm_interconnect_0:game_cpu_data_master_waitrequest -> game_cpu:d_waitrequest
	wire         game_cpu_data_master_debugaccess;                          // game_cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:game_cpu_data_master_debugaccess
	wire  [28:0] game_cpu_data_master_address;                              // game_cpu:d_address -> mm_interconnect_0:game_cpu_data_master_address
	wire   [3:0] game_cpu_data_master_byteenable;                           // game_cpu:d_byteenable -> mm_interconnect_0:game_cpu_data_master_byteenable
	wire         game_cpu_data_master_read;                                 // game_cpu:d_read -> mm_interconnect_0:game_cpu_data_master_read
	wire         game_cpu_data_master_write;                                // game_cpu:d_write -> mm_interconnect_0:game_cpu_data_master_write
	wire  [31:0] game_cpu_data_master_writedata;                            // game_cpu:d_writedata -> mm_interconnect_0:game_cpu_data_master_writedata
	wire  [31:0] game_cpu_instruction_master_readdata;                      // mm_interconnect_0:game_cpu_instruction_master_readdata -> game_cpu:i_readdata
	wire         game_cpu_instruction_master_waitrequest;                   // mm_interconnect_0:game_cpu_instruction_master_waitrequest -> game_cpu:i_waitrequest
	wire  [28:0] game_cpu_instruction_master_address;                       // game_cpu:i_address -> mm_interconnect_0:game_cpu_instruction_master_address
	wire         game_cpu_instruction_master_read;                          // game_cpu:i_read -> mm_interconnect_0:game_cpu_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_avalon_game_interface_avl_chipselect;    // mm_interconnect_0:avalon_game_interface_avl_chipselect -> avalon_game_interface:AVL_CS
	wire  [31:0] mm_interconnect_0_avalon_game_interface_avl_readdata;      // avalon_game_interface:AVL_READDATA -> mm_interconnect_0:avalon_game_interface_avl_readdata
	wire   [5:0] mm_interconnect_0_avalon_game_interface_avl_address;       // mm_interconnect_0:avalon_game_interface_avl_address -> avalon_game_interface:AVL_ADDR
	wire         mm_interconnect_0_avalon_game_interface_avl_read;          // mm_interconnect_0:avalon_game_interface_avl_read -> avalon_game_interface:AVL_READ
	wire   [3:0] mm_interconnect_0_avalon_game_interface_avl_byteenable;    // mm_interconnect_0:avalon_game_interface_avl_byteenable -> avalon_game_interface:AVL_BYTE_EN
	wire         mm_interconnect_0_avalon_game_interface_avl_write;         // mm_interconnect_0:avalon_game_interface_avl_write -> avalon_game_interface:AVL_WRITE
	wire  [31:0] mm_interconnect_0_avalon_game_interface_avl_writedata;     // mm_interconnect_0:avalon_game_interface_avl_writedata -> avalon_game_interface:AVL_WRITEDATA
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;       // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;        // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_game_cpu_debug_mem_slave_readdata;       // game_cpu:debug_mem_slave_readdata -> mm_interconnect_0:game_cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_game_cpu_debug_mem_slave_waitrequest;    // game_cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:game_cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_game_cpu_debug_mem_slave_debugaccess;    // mm_interconnect_0:game_cpu_debug_mem_slave_debugaccess -> game_cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_game_cpu_debug_mem_slave_address;        // mm_interconnect_0:game_cpu_debug_mem_slave_address -> game_cpu:debug_mem_slave_address
	wire         mm_interconnect_0_game_cpu_debug_mem_slave_read;           // mm_interconnect_0:game_cpu_debug_mem_slave_read -> game_cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_game_cpu_debug_mem_slave_byteenable;     // mm_interconnect_0:game_cpu_debug_mem_slave_byteenable -> game_cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_game_cpu_debug_mem_slave_write;          // mm_interconnect_0:game_cpu_debug_mem_slave_write -> game_cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_game_cpu_debug_mem_slave_writedata;      // mm_interconnect_0:game_cpu_debug_mem_slave_writedata -> game_cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_system_pll_pll_slave_readdata;           // system_pll:readdata -> mm_interconnect_0:system_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_system_pll_pll_slave_address;            // mm_interconnect_0:system_pll_pll_slave_address -> system_pll:address
	wire         mm_interconnect_0_system_pll_pll_slave_read;               // mm_interconnect_0:system_pll_pll_slave_read -> system_pll:read
	wire         mm_interconnect_0_system_pll_pll_slave_write;              // mm_interconnect_0:system_pll_pll_slave_write -> system_pll:write
	wire  [31:0] mm_interconnect_0_system_pll_pll_slave_writedata;          // mm_interconnect_0:system_pll_pll_slave_writedata -> system_pll:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                     // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                       // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                    // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                        // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                           // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                     // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                  // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                          // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                      // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_otg_hpi_address_s1_chipselect;           // mm_interconnect_0:otg_hpi_address_s1_chipselect -> otg_hpi_address:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_address_s1_readdata;             // otg_hpi_address:readdata -> mm_interconnect_0:otg_hpi_address_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_address_s1_address;              // mm_interconnect_0:otg_hpi_address_s1_address -> otg_hpi_address:address
	wire         mm_interconnect_0_otg_hpi_address_s1_write;                // mm_interconnect_0:otg_hpi_address_s1_write -> otg_hpi_address:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_address_s1_writedata;            // mm_interconnect_0:otg_hpi_address_s1_writedata -> otg_hpi_address:writedata
	wire         mm_interconnect_0_otg_hpi_data_s1_chipselect;              // mm_interconnect_0:otg_hpi_data_s1_chipselect -> otg_hpi_data:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_data_s1_readdata;                // otg_hpi_data:readdata -> mm_interconnect_0:otg_hpi_data_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_data_s1_address;                 // mm_interconnect_0:otg_hpi_data_s1_address -> otg_hpi_data:address
	wire         mm_interconnect_0_otg_hpi_data_s1_write;                   // mm_interconnect_0:otg_hpi_data_s1_write -> otg_hpi_data:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_data_s1_writedata;               // mm_interconnect_0:otg_hpi_data_s1_writedata -> otg_hpi_data:writedata
	wire         mm_interconnect_0_otg_hpi_r_s1_chipselect;                 // mm_interconnect_0:otg_hpi_r_s1_chipselect -> otg_hpi_r:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_r_s1_readdata;                   // otg_hpi_r:readdata -> mm_interconnect_0:otg_hpi_r_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_r_s1_address;                    // mm_interconnect_0:otg_hpi_r_s1_address -> otg_hpi_r:address
	wire         mm_interconnect_0_otg_hpi_r_s1_write;                      // mm_interconnect_0:otg_hpi_r_s1_write -> otg_hpi_r:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_r_s1_writedata;                  // mm_interconnect_0:otg_hpi_r_s1_writedata -> otg_hpi_r:writedata
	wire         mm_interconnect_0_otg_hpi_w_s1_chipselect;                 // mm_interconnect_0:otg_hpi_w_s1_chipselect -> otg_hpi_w:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_w_s1_readdata;                   // otg_hpi_w:readdata -> mm_interconnect_0:otg_hpi_w_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_w_s1_address;                    // mm_interconnect_0:otg_hpi_w_s1_address -> otg_hpi_w:address
	wire         mm_interconnect_0_otg_hpi_w_s1_write;                      // mm_interconnect_0:otg_hpi_w_s1_write -> otg_hpi_w:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_w_s1_writedata;                  // mm_interconnect_0:otg_hpi_w_s1_writedata -> otg_hpi_w:writedata
	wire         mm_interconnect_0_otg_hpi_cs_s1_chipselect;                // mm_interconnect_0:otg_hpi_cs_s1_chipselect -> otg_hpi_cs:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_cs_s1_readdata;                  // otg_hpi_cs:readdata -> mm_interconnect_0:otg_hpi_cs_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_cs_s1_address;                   // mm_interconnect_0:otg_hpi_cs_s1_address -> otg_hpi_cs:address
	wire         mm_interconnect_0_otg_hpi_cs_s1_write;                     // mm_interconnect_0:otg_hpi_cs_s1_write -> otg_hpi_cs:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_cs_s1_writedata;                 // mm_interconnect_0:otg_hpi_cs_s1_writedata -> otg_hpi_cs:writedata
	wire         mm_interconnect_0_otg_hpi_reset_s1_chipselect;             // mm_interconnect_0:otg_hpi_reset_s1_chipselect -> otg_hpi_reset:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_reset_s1_readdata;               // otg_hpi_reset:readdata -> mm_interconnect_0:otg_hpi_reset_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_reset_s1_address;                // mm_interconnect_0:otg_hpi_reset_s1_address -> otg_hpi_reset:address
	wire         mm_interconnect_0_otg_hpi_reset_s1_write;                  // mm_interconnect_0:otg_hpi_reset_s1_write -> otg_hpi_reset:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_reset_s1_writedata;              // mm_interconnect_0:otg_hpi_reset_s1_writedata -> otg_hpi_reset:writedata
	wire  [31:0] mm_interconnect_0_frame_sync_s1_readdata;                  // frame_sync:readdata -> mm_interconnect_0:frame_sync_s1_readdata
	wire   [1:0] mm_interconnect_0_frame_sync_s1_address;                   // mm_interconnect_0:frame_sync_s1_address -> frame_sync:address
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] game_cpu_irq_irq;                                          // irq_mapper:sender_irq -> game_cpu:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [avalon_game_interface:RESET, frame_sync:reset_n, jtag_uart:rst_n, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, otg_hpi_address:reset_n, otg_hpi_cs:reset_n, otg_hpi_data:reset_n, otg_hpi_r:reset_n, otg_hpi_reset:reset_n, otg_hpi_w:reset_n, sysid_qsys:reset_n, system_pll:reset]
	wire         game_cpu_debug_reset_request_reset;                        // game_cpu:debug_reset_request -> [rst_controller:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [game_cpu:reset_n, irq_mapper:reset, mm_interconnect_0:game_cpu_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset_req;                    // rst_controller_001:reset_req -> [game_cpu:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> [mm_interconnect_0:sdram_reset_reset_bridge_in_reset_reset, sdram:reset_n]

	avalon_game_interface avalon_game_interface (
		.CLK           (clk_clk),                                                //  clock.clk
		.RESET         (rst_controller_reset_out_reset),                         //  reset.reset
		.AVL_READ      (mm_interconnect_0_avalon_game_interface_avl_read),       //    avl.read
		.AVL_WRITE     (mm_interconnect_0_avalon_game_interface_avl_write),      //       .write
		.AVL_WRITEDATA (mm_interconnect_0_avalon_game_interface_avl_writedata),  //       .writedata
		.AVL_READDATA  (mm_interconnect_0_avalon_game_interface_avl_readdata),   //       .readdata
		.AVL_ADDR      (mm_interconnect_0_avalon_game_interface_avl_address),    //       .address
		.AVL_BYTE_EN   (mm_interconnect_0_avalon_game_interface_avl_byteenable), //       .byteenable
		.AVL_CS        (mm_interconnect_0_avalon_game_interface_avl_chipselect), //       .chipselect
		.EXPORT_DATA   (gamefile_export_data)                                    // EXPORT.export_data
	);

	final_soc_frame_sync frame_sync (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_frame_sync_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_frame_sync_s1_readdata), //                    .readdata
		.in_port  (frame_sync_export)                         // external_connection.export
	);

	final_soc_game_cpu game_cpu (
		.clk                                 (clk_clk),                                                //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (game_cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (game_cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (game_cpu_data_master_read),                              //                          .read
		.d_readdata                          (game_cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (game_cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (game_cpu_data_master_write),                             //                          .write
		.d_writedata                         (game_cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (game_cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (game_cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (game_cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (game_cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (game_cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (game_cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (game_cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_game_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_game_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_game_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_game_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_game_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_game_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_game_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_game_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                        // custom_instruction_master.readra
	);

	final_soc_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	final_soc_otg_hpi_address otg_hpi_address (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_address_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_address_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_address_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_address_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_address_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_address_export)                           // external_connection.export
	);

	final_soc_otg_hpi_cs otg_hpi_cs (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_cs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_cs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_cs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_cs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_cs_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_cs_export)                           // external_connection.export
	);

	final_soc_otg_hpi_data otg_hpi_data (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_data_s1_readdata),   //                    .readdata
		.in_port    (otg_hpi_data_in_port),                         // external_connection.export
		.out_port   (otg_hpi_data_out_port)                         //                    .export
	);

	final_soc_otg_hpi_cs otg_hpi_r (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_r_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_r_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_r_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_r_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_r_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_r_export)                           // external_connection.export
	);

	final_soc_otg_hpi_cs otg_hpi_reset (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_reset_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_reset_export)                           // external_connection.export
	);

	final_soc_otg_hpi_cs otg_hpi_w (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_w_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_w_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_w_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_w_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_w_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_w_export)                           // external_connection.export
	);

	final_soc_sdram sdram (
		.clk            (system_pll_c0_clk),                        //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	final_soc_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	final_soc_system_pll system_pll (
		.clk                (clk_clk),                                          //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                   // inclk_interface_reset.reset
		.read               (mm_interconnect_0_system_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_system_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_system_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_system_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_system_pll_pll_slave_writedata), //                      .writedata
		.c0                 (system_pll_c0_clk),                                //                    c0.clk
		.c1                 (sdram_clk_clk),                                    //                    c1.clk
		.scandone           (),                                                 //           (terminated)
		.scandataout        (),                                                 //           (terminated)
		.areset             (1'b0),                                             //           (terminated)
		.locked             (),                                                 //           (terminated)
		.phasedone          (),                                                 //           (terminated)
		.phasecounterselect (4'b0000),                                          //           (terminated)
		.phaseupdown        (1'b0),                                             //           (terminated)
		.phasestep          (1'b0),                                             //           (terminated)
		.scanclk            (1'b0),                                             //           (terminated)
		.scanclkena         (1'b0),                                             //           (terminated)
		.scandata           (1'b0),                                             //           (terminated)
		.configupdate       (1'b0)                                              //           (terminated)
	);

	final_soc_mm_interconnect_0 mm_interconnect_0 (
		.system_clk_clk_clk                          (clk_clk),                                                   //                        system_clk_clk.clk
		.system_pll_c0_clk                           (system_pll_c0_clk),                                         //                         system_pll_c0.clk
		.game_cpu_reset_reset_bridge_in_reset_reset  (rst_controller_001_reset_out_reset),                        //  game_cpu_reset_reset_bridge_in_reset.reset
		.jtag_uart_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // jtag_uart_reset_reset_bridge_in_reset.reset
		.sdram_reset_reset_bridge_in_reset_reset     (rst_controller_002_reset_out_reset),                        //     sdram_reset_reset_bridge_in_reset.reset
		.game_cpu_data_master_address                (game_cpu_data_master_address),                              //                  game_cpu_data_master.address
		.game_cpu_data_master_waitrequest            (game_cpu_data_master_waitrequest),                          //                                      .waitrequest
		.game_cpu_data_master_byteenable             (game_cpu_data_master_byteenable),                           //                                      .byteenable
		.game_cpu_data_master_read                   (game_cpu_data_master_read),                                 //                                      .read
		.game_cpu_data_master_readdata               (game_cpu_data_master_readdata),                             //                                      .readdata
		.game_cpu_data_master_write                  (game_cpu_data_master_write),                                //                                      .write
		.game_cpu_data_master_writedata              (game_cpu_data_master_writedata),                            //                                      .writedata
		.game_cpu_data_master_debugaccess            (game_cpu_data_master_debugaccess),                          //                                      .debugaccess
		.game_cpu_instruction_master_address         (game_cpu_instruction_master_address),                       //           game_cpu_instruction_master.address
		.game_cpu_instruction_master_waitrequest     (game_cpu_instruction_master_waitrequest),                   //                                      .waitrequest
		.game_cpu_instruction_master_read            (game_cpu_instruction_master_read),                          //                                      .read
		.game_cpu_instruction_master_readdata        (game_cpu_instruction_master_readdata),                      //                                      .readdata
		.avalon_game_interface_avl_address           (mm_interconnect_0_avalon_game_interface_avl_address),       //             avalon_game_interface_avl.address
		.avalon_game_interface_avl_write             (mm_interconnect_0_avalon_game_interface_avl_write),         //                                      .write
		.avalon_game_interface_avl_read              (mm_interconnect_0_avalon_game_interface_avl_read),          //                                      .read
		.avalon_game_interface_avl_readdata          (mm_interconnect_0_avalon_game_interface_avl_readdata),      //                                      .readdata
		.avalon_game_interface_avl_writedata         (mm_interconnect_0_avalon_game_interface_avl_writedata),     //                                      .writedata
		.avalon_game_interface_avl_byteenable        (mm_interconnect_0_avalon_game_interface_avl_byteenable),    //                                      .byteenable
		.avalon_game_interface_avl_chipselect        (mm_interconnect_0_avalon_game_interface_avl_chipselect),    //                                      .chipselect
		.frame_sync_s1_address                       (mm_interconnect_0_frame_sync_s1_address),                   //                         frame_sync_s1.address
		.frame_sync_s1_readdata                      (mm_interconnect_0_frame_sync_s1_readdata),                  //                                      .readdata
		.game_cpu_debug_mem_slave_address            (mm_interconnect_0_game_cpu_debug_mem_slave_address),        //              game_cpu_debug_mem_slave.address
		.game_cpu_debug_mem_slave_write              (mm_interconnect_0_game_cpu_debug_mem_slave_write),          //                                      .write
		.game_cpu_debug_mem_slave_read               (mm_interconnect_0_game_cpu_debug_mem_slave_read),           //                                      .read
		.game_cpu_debug_mem_slave_readdata           (mm_interconnect_0_game_cpu_debug_mem_slave_readdata),       //                                      .readdata
		.game_cpu_debug_mem_slave_writedata          (mm_interconnect_0_game_cpu_debug_mem_slave_writedata),      //                                      .writedata
		.game_cpu_debug_mem_slave_byteenable         (mm_interconnect_0_game_cpu_debug_mem_slave_byteenable),     //                                      .byteenable
		.game_cpu_debug_mem_slave_waitrequest        (mm_interconnect_0_game_cpu_debug_mem_slave_waitrequest),    //                                      .waitrequest
		.game_cpu_debug_mem_slave_debugaccess        (mm_interconnect_0_game_cpu_debug_mem_slave_debugaccess),    //                                      .debugaccess
		.jtag_uart_avalon_jtag_slave_address         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //           jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                      .write
		.jtag_uart_avalon_jtag_slave_read            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                      .read
		.jtag_uart_avalon_jtag_slave_readdata        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                      .readdata
		.jtag_uart_avalon_jtag_slave_writedata       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                      .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                      .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                      .chipselect
		.otg_hpi_address_s1_address                  (mm_interconnect_0_otg_hpi_address_s1_address),              //                    otg_hpi_address_s1.address
		.otg_hpi_address_s1_write                    (mm_interconnect_0_otg_hpi_address_s1_write),                //                                      .write
		.otg_hpi_address_s1_readdata                 (mm_interconnect_0_otg_hpi_address_s1_readdata),             //                                      .readdata
		.otg_hpi_address_s1_writedata                (mm_interconnect_0_otg_hpi_address_s1_writedata),            //                                      .writedata
		.otg_hpi_address_s1_chipselect               (mm_interconnect_0_otg_hpi_address_s1_chipselect),           //                                      .chipselect
		.otg_hpi_cs_s1_address                       (mm_interconnect_0_otg_hpi_cs_s1_address),                   //                         otg_hpi_cs_s1.address
		.otg_hpi_cs_s1_write                         (mm_interconnect_0_otg_hpi_cs_s1_write),                     //                                      .write
		.otg_hpi_cs_s1_readdata                      (mm_interconnect_0_otg_hpi_cs_s1_readdata),                  //                                      .readdata
		.otg_hpi_cs_s1_writedata                     (mm_interconnect_0_otg_hpi_cs_s1_writedata),                 //                                      .writedata
		.otg_hpi_cs_s1_chipselect                    (mm_interconnect_0_otg_hpi_cs_s1_chipselect),                //                                      .chipselect
		.otg_hpi_data_s1_address                     (mm_interconnect_0_otg_hpi_data_s1_address),                 //                       otg_hpi_data_s1.address
		.otg_hpi_data_s1_write                       (mm_interconnect_0_otg_hpi_data_s1_write),                   //                                      .write
		.otg_hpi_data_s1_readdata                    (mm_interconnect_0_otg_hpi_data_s1_readdata),                //                                      .readdata
		.otg_hpi_data_s1_writedata                   (mm_interconnect_0_otg_hpi_data_s1_writedata),               //                                      .writedata
		.otg_hpi_data_s1_chipselect                  (mm_interconnect_0_otg_hpi_data_s1_chipselect),              //                                      .chipselect
		.otg_hpi_r_s1_address                        (mm_interconnect_0_otg_hpi_r_s1_address),                    //                          otg_hpi_r_s1.address
		.otg_hpi_r_s1_write                          (mm_interconnect_0_otg_hpi_r_s1_write),                      //                                      .write
		.otg_hpi_r_s1_readdata                       (mm_interconnect_0_otg_hpi_r_s1_readdata),                   //                                      .readdata
		.otg_hpi_r_s1_writedata                      (mm_interconnect_0_otg_hpi_r_s1_writedata),                  //                                      .writedata
		.otg_hpi_r_s1_chipselect                     (mm_interconnect_0_otg_hpi_r_s1_chipselect),                 //                                      .chipselect
		.otg_hpi_reset_s1_address                    (mm_interconnect_0_otg_hpi_reset_s1_address),                //                      otg_hpi_reset_s1.address
		.otg_hpi_reset_s1_write                      (mm_interconnect_0_otg_hpi_reset_s1_write),                  //                                      .write
		.otg_hpi_reset_s1_readdata                   (mm_interconnect_0_otg_hpi_reset_s1_readdata),               //                                      .readdata
		.otg_hpi_reset_s1_writedata                  (mm_interconnect_0_otg_hpi_reset_s1_writedata),              //                                      .writedata
		.otg_hpi_reset_s1_chipselect                 (mm_interconnect_0_otg_hpi_reset_s1_chipselect),             //                                      .chipselect
		.otg_hpi_w_s1_address                        (mm_interconnect_0_otg_hpi_w_s1_address),                    //                          otg_hpi_w_s1.address
		.otg_hpi_w_s1_write                          (mm_interconnect_0_otg_hpi_w_s1_write),                      //                                      .write
		.otg_hpi_w_s1_readdata                       (mm_interconnect_0_otg_hpi_w_s1_readdata),                   //                                      .readdata
		.otg_hpi_w_s1_writedata                      (mm_interconnect_0_otg_hpi_w_s1_writedata),                  //                                      .writedata
		.otg_hpi_w_s1_chipselect                     (mm_interconnect_0_otg_hpi_w_s1_chipselect),                 //                                      .chipselect
		.sdram_s1_address                            (mm_interconnect_0_sdram_s1_address),                        //                              sdram_s1.address
		.sdram_s1_write                              (mm_interconnect_0_sdram_s1_write),                          //                                      .write
		.sdram_s1_read                               (mm_interconnect_0_sdram_s1_read),                           //                                      .read
		.sdram_s1_readdata                           (mm_interconnect_0_sdram_s1_readdata),                       //                                      .readdata
		.sdram_s1_writedata                          (mm_interconnect_0_sdram_s1_writedata),                      //                                      .writedata
		.sdram_s1_byteenable                         (mm_interconnect_0_sdram_s1_byteenable),                     //                                      .byteenable
		.sdram_s1_readdatavalid                      (mm_interconnect_0_sdram_s1_readdatavalid),                  //                                      .readdatavalid
		.sdram_s1_waitrequest                        (mm_interconnect_0_sdram_s1_waitrequest),                    //                                      .waitrequest
		.sdram_s1_chipselect                         (mm_interconnect_0_sdram_s1_chipselect),                     //                                      .chipselect
		.sysid_qsys_control_slave_address            (mm_interconnect_0_sysid_qsys_control_slave_address),        //              sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata           (mm_interconnect_0_sysid_qsys_control_slave_readdata),       //                                      .readdata
		.system_pll_pll_slave_address                (mm_interconnect_0_system_pll_pll_slave_address),            //                  system_pll_pll_slave.address
		.system_pll_pll_slave_write                  (mm_interconnect_0_system_pll_pll_slave_write),              //                                      .write
		.system_pll_pll_slave_read                   (mm_interconnect_0_system_pll_pll_slave_read),               //                                      .read
		.system_pll_pll_slave_readdata               (mm_interconnect_0_system_pll_pll_slave_readdata),           //                                      .readdata
		.system_pll_pll_slave_writedata              (mm_interconnect_0_system_pll_pll_slave_writedata)           //                                      .writedata
	);

	final_soc_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (game_cpu_irq_irq)                    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (game_cpu_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (game_cpu_debug_reset_request_reset), // reset_in1.reset
		.clk            (system_pll_c0_clk),                  //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
